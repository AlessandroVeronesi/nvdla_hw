`ifndef __COMMONS_VH__
`define __COMMONS_VH__

`define FIFOGEN_MASTER_CLK_GATING_DISABLED
`define SYNTHESIS
`define FPGA
`define NV_FPGA_FIGOGEN
`define VLIB_BYPASS_POWER_CG

`endif